b0VIM 8.0      N�cB �l  root                                    fraude.omegasin.ma                      /var/www/veopro/VEO/views.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp(           �                            b       �                     S       �                     d       9                    d       �                    a                            a       b             !       _       �             "       ]       "             #       Y                    $       ]       �             %       \       5             &       V       �             '       [       �             (       O       B                    O       �             )       d       �                    n       D                    v       �                    Z       (                    `       �             	       U       �             
       _       7                    a       �                    ^       �                    [       U	                    [       �	                    [       
                    X       f
                    [       �
                    Z                           U       s                    V       �                    Y                           K       w                    U       �                    x                           w       �                    h                           -       n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     >     �       �  �  h  .    �  �  �  r  f  e  *  )  (  '  &    �  �  z  y  `  J    �  �  �  �  O    �  �  �  k  O  G      �
  �
  �
  �
  �
  �
  �
  u
  S
  3
  
  
  �	  �	  �	  �	  �	  �	  }	  ^	  @	  /	  	  	  	  	  �  �  �  �  �  p  o  8  '  �  �  �  �  c  C  5           �  �  �  P    	  �  �  �  �  �  �  {  c  O  ;      �  �  �  �  v  ^  5      �  �  �  �  �  u  d  Z  A  1  0  /      �  w  s  `  H  >  =                            NBD=0     list_Veo_recente=[]     NBDAT=nbrDAT()         Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def inis(request): @login_required       return stri         stri=float(stri)     else:         stri=0.0     if stri == "" or stri == "'0.0'" or stri  == None: def str_to_float(stri): #Convertir Rate fraude de string to float               return a             a=test(a)             a=add_zero(a)         if (a != '' and not(a is None)):         a=remove_WW0(a)         a=remove_WW(a)         a=remove_zerostart(a)         a=a.replace('-','')         a=a.replace(".", "")         a=a.replace("'", "")         a=a.replace("/", "")         a=a.replace(" ", "")         a=a.upper()         a=a.strip()         a=remove_EAD(a)     if a!=None: def Preprocessing_Imm (a): #Preprocessing "Immatriculation" (Appeler toutes les fcts défénies)           return a     else:         return ""     if ((len(b) == len(a)) or ((len(c) == len(a)))):     c=''.join(i for i in a if not (i.isdigit()))     b=''.join(i for i in a if i.isdigit()) def test(a): #Enlever les imm qui contient que des chiffres ou bien que des caractères          return a     else:             return a         else:             return ''.join(res)             res.append(a[-1])             res.append("0")             res=list(a)[0:-1]         if (a[-1].isdigit() and (not a[-2].isdigit())):     if (len(a) <= 2 or a != '' or not (a is None)): def add_zero(a): #Ajouter le le zéro après le caractère (B7 ==> B07)          return a     else:         return ''.join(list(a)[3:])     if (a.startswith("EAD")): def remove_EAD(a): #Enlever le mot "EAD" s'il existe          return a     else:         return a         a="WW"+a         a=remove_zerostart(a)         a=''.join(list(a)[2:])     if a.startswith("WW0"): def remove_WW0(a): #Enlever les zeros après les "WW" de début          return a     else:             return "WW"+a         else :             return a         if(a.startswith("WW")):         a= ''.join(list(a)[0:-2])     if a.endswith("WW"): def remove_WW(a): #Enlever les "WW" à la fin      return val         val = ''.join(l)         i=i+1         l[0]=''         l=list(val)     while (val.startswith('0') and i<len(val)):     i=0 def remove_zerostart (val): #Enlever les zéros de début ################################################################### Nettoyage des immatriculations          return (dtV - dtE).days         dtV = datetime.strptime(dtV, "%d %b, %Y %H:%M:%S").date()         dtE = datetime.strptime(dtE, "%d/%m/%Y").date()     if (dtV and dtE): def inter_dt2(dtV , dtE):         return abs(dtV - dtE).days         dtE = datetime.strptime(dtE, "%d/%m/%Y").date()         dtV = datetime.strptime(dtV, "%d/%m/%Y").date()     if (dtV and dtE): def inter_dt(dtV , dtE):      return a     a=a.replace(' ','').replace('-','').replace('_','').replace(',','').replace('.','').replace('*','') def net_numch(a): # nettoyage  de  numéro de  chassis     from django.core.serializers.json import DjangoJSONEncoder  import json from django.core.serializers import serialize from django.http import HttpResponse from django.core.paginator import Paginator import datetime from django.http import HttpResponseRedirect from django.contrib.auth.decorators import login_required from .models import Veodata, Assistance, Bris_De_Glace, Veoservices,veotest from django.shortcuts import render, get_object_or_404 from os import lseek ad  �  �     -       �  �  �  �  �  y  o  c  [  Z    �  �  �  �  b  ?  �  �  g  [  P  :  #  n  [  T  *    �  I  +    _
  J
  -
  
  �	  �	  S	  ;	  1	  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         return HttpResponse(response, content_type='text/json')     response = jsls         response = json.dumps([{'Error':'Invalid Token'}])"""     else:         response = jsls     """if 'authorization' in request.headers and request.headers['authorization'] == 'Basic VeosmartAyODkwNUUteWx1LTIwTEM5RzRNQFZFT1NNQVJUV0FGQQ==':          #jsl = [line for line in jsls]     #jsls = json.loads(jsls)     #jsls = json.dumps(jsls)     jsls.append(']')     jsls.append({'Dossier':l.Dossier,'Pourcentage Fraude':l.RateFraude,'Procédure':l.Procédure,'Statut':l.Statut,'Date Création':l.Date_création,'Statut doute':l.statutdoute})      jsls.append(",")               jsls.append(js)               js={'Dossier':j.Dossier,'Pourcentage Fraude':j.RateFraude,'Procédure':j.Procédure,'Statut':j.Statut,'Date Création':j.Date_création,'Statut doute':j.statutdoute}             jsls.append(",")             N=N+1         if  j != k and j != l and N<1001:            for j  in  ls:     jsls.append({'Dossier':k.Dossier,'Pourcentage Fraude':k.RateFraude,'Procédure':k.Procédure,'Statut':k.Statut,'Date Création':k.Date_création,'Statut doute':k.statutdoute})      jsls.append('[')       l=ls[len(ls)-1]                  k=ls[0]                 ls.append(i)             if ((Today_DateVeo-Date_création).days<=15) and i.RateFraude not in [0,'0.0',None]:             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_Veoservices:     Rate=0     list_Veoservices=Veoservices.objects.all()     NBD=0     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')      N=2     jsls=[]     ls=[]     veoservice=Veoservices.objects.all()      def get_dossiers(request):       return HttpResponse(response, content_type='text/json') ad     m     O       �  l  N  &  �  �  q  X  =  $    �  �  �  Z      �  �  i  ;    �
  �
  �
  �
  �
  �
  e
  @
  �	  �	  �	  �	  	  �  �  �  �  �  �  m  N  %    g  1  
  	  �  �  u  P  O  8    �  �  �  \  6    �  \  L  /      �  �  �  �  q  ,    �  �  �  m  g                                   i.RateFraude = str_to_float(i.RateFraude)         if (i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) :              for i in list_Veoservices:             list_inst.append(i)         if i.Statut =="Dossier en instruction" and "D" in i.Dossier:     for i in list_Veoservicesall:     list_Veoservicesall= Veoservices.objects.all()     list_Veoservices=DosAff()     list_inst=[]     list_Veo_recente=[]     NBDT=nbrDT()     NBD=nbrDAT() def dossiersAtrait(request): @login_required     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT}    # veoD = paginator.get_page(pageD)    # pageD = request.GET.get('pageD')    # paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]      veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)              list_Veo_recente.append(i)             i.RateFraude = str_to_float(i.RateFraude)         if (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté") and i.Statut!="Changement de procédure" and  i.Statut!="Dossier sans suite" :     for i in list_Veoservices:     Veoservice=Veoservices.objects.all()     list_Veoservices=DosTAff()     list_Veo_recente=[]     NBDT=nbrDT()     NBD=nbrDAT() def dossierstrait(request): @login_required      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()           veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                         i.RateFraude=str_to_float(i.RateFraude)                         list_Veo_recente.append(i)                     if (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté") and i.Statut!="Changement de procédure" and  i.Statut!="Dossier sans suite" and i.RateFraude not in [0,'0.0',None,'5.0','10.0'] and i not in list_Veo_recente:                 if ((Today_DateVeo-Date_création).days<=100):                 Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')             if i.Date_création!=None:         for i in liste:             liste=liste1+liste2         else:             liste=liste1         elif liste2==None:             liste=liste2         if liste1==None:         liste1=list(Veoservices.objects.filter(Immatriculation__icontains=query))         liste2=list(Veoservices.objects.filter(Dossier__icontains=query))         query=request.GET.get('search')     if request.method=='GET':     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') ad     �     n       �  �  �  �  �  �  �  �  v  Z  G  '  �  �  �  �  y  Y  C  #  �  �  �  �  �  l  L  6    �
  �
  �
  �
  h
  H
  2
  
  �	  �	  �	  �	  d	  D	  .	  	  �  �  �  �  ]  =  &    �  �  �  �  S  3  .    �  �  �  �  q  Q    �  �  �  �  �  ~  ^  Y  T  1    �  �  }  N  M  L  K  J  I  D  )      �  �  �  �    _  I  )  �  �  �  �  {  [  R  <    �  �                                          if i.R4 != None and i.R4 != "":         for i in listedossiers:     elif (ch =="R4"):                          liste.append(i)             if i.R3 != None and i.R3 != "":         for i in listedossiers:     elif (ch =="R3"):                 liste.append(i)             if i.R2 != None and i.R2 != "":         for i in listedossiers:     elif (ch =="R2"):                 liste.append(i)             if i.R1 != None and i.R1 != "":         for i in listedossiers:     if (ch=="R1"):     listedossiers =DosAT()     liste=[]          ch=request.GET.get('reg') def filtre_regAT(request):               return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDossiers":NBDAT,"list_Veo_recente": veopg }     NBDAT=nbrDAT()         veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(liste,9)                           liste.append(i)             if i.R14 != None and i.R14 != "":         for i in listedossiers:     elif (ch =="R14"):                                   liste.append(i)             if i.R13 != None and "doute rejeté" in i.R13 :         for i in listedossiers:     elif (ch =="R13_rejete"):                  liste.append(i)             if i.R13 != None and "doute confirmé" in i.R13 :         for i in listedossiers:     elif (ch =="R13_confirme"):                      liste.append(i)             if i.R12 != None and i.R12 != "":         for i in listedossiers:     elif (ch =="R12"):                 liste.append(i)             if i.R11 != None and i.R11 != "":         for i in listedossiers:     elif (ch =="R11"):                 liste.append(i)             if i.R10 != None and i.R10 != "":         for i in listedossiers:     elif (ch =="R10"):                 liste.append(i)             if i.R9 != None and i.R9 != "":         for i in listedossiers:     elif (ch =="R9"):                 liste.append(i)             if i.R8 != None and i.R8 != "":         for i in listedossiers:     elif (ch =="R8"):                 liste.append(i)             if i.R7 != None and i.R7 != "":         for i in listedossiers:     elif (ch =="R7"):                 liste.append(i)             if i.R6 != None and i.R6 != "":         for i in listedossiers:     elif (ch =="R6"):                 liste.append(i)             if i.R5 != None and i.R5 != "":         for i in listedossiers:     elif (ch =="R5"):                 liste.append(i)             if i.R4 != None and i.R4 != "":         for i in listedossiers:     elif (ch =="R4"):                          liste.append(i)             if i.R3 != None and i.R3 != "":         for i in listedossiers:     elif (ch =="R3"):                 liste.append(i)             if i.R2 != None and i.R2 != "":         for i in listedossiers:     elif (ch =="R2"):                 liste.append(i)             if i.R1 != None and i.R1 != "":         for i in listedossiers:     if (ch=="R1"):     listedossiers =DosAff()     liste=[]          ch=request.GET.get('reg') def filtre_reg(request):            return render(request,"detail.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"Veo":Veo,"Rate":Rate ,"R1": R1,"R1_P": R1_P, "R1_A":R1_A, "R2":R2, "R2_DDA":R2_DDA, "R2_DS":R2_DS,"R3":R3, "R3_DDA":R3_DDA, "R3_DS":R3_DS, "R4":R4, "R4_SP":R4_SP, "R4_SA":R4_SA,"R5":R5 ,"R5_Assis":R5_Assis ,"R6":R6,"R6_Assis1":R6_Assis1 ,"R6_Assis2":R6_Assis2,"R7":R7,"R7_P":R7_P,"R7_A":R7_A, "R9_DFP":R9_DFP, "R9_DS":R9_DS, "R9":R9,"R8":R8,"NBDossiers":NBD,"R11":R11, "R10_Dos":R10_Dos,"R10":R10 , "R12_Dos":R12_Dos,"R12":R12 , "R14":R14, "R13_Dos":R13_Dos,"R13":R13 } ad          v       �  �  �  ~  ^  H  (  �  �  �  �  z  Z  D  $  �  �  �  �  v  V  ?    �  �  �  �  l  L  5    �  �  �  �  �  F  &  %    �
  �
  �
  �
  y
  b
  B
  
  �	  �	  �	  �	  �	  s	  n	  	  	  �  �  �  �  �  �  �  �  q  ^  >    �  �  �  �  p  Z  :    �  �  �  �  �  c  M  -    �  �  �    _  I  )  �  �  �  �  {  [  E  %  �  �  �  �  t  T  =    �  �  �  �  j  J  G  '                                 for i in listedossiers:     elif (ch =="R13_confirme"):                    liste.append(i)             if i.R12 != None and i.R12 != "":         for i in listedossiers:     elif (ch =="R12"):                 liste.append(i)             if i.R11 != None and i.R11 != "":         for i in listedossiers:     elif (ch =="R11"):                 liste.append(i)             if i.R10 != None and i.R10 != "":         for i in listedossiers:     elif (ch =="R10"):                 liste.append(i)             if i.R9 != None and i.R9 != "":         for i in listedossiers:     elif (ch =="R9"):                 liste.append(i)             if i.R8 != None and i.R8 != "":         for i in listedossiers:     elif (ch =="R8"):                 liste.append(i)             if i.R7 != None and i.R7 != "":         for i in listedossiers:     elif (ch =="R7"):                 liste.append(i)             if i.R6 != None and i.R6 != "":         for i in listedossiers:     elif (ch =="R6"):                 liste.append(i)             if i.R5 != None and i.R5 != "":         for i in listedossiers:     elif (ch =="R5"):                 liste.append(i)             if i.R4 != None and i.R4 != "":         for i in listedossiers:     elif (ch =="R4"):                          liste.append(i)             if i.R3 != None and i.R3 != "":         for i in listedossiers:     elif (ch =="R3"):                 liste.append(i)             if i.R2 != None and i.R2 != "":         for i in listedossiers:     elif (ch =="R2"):                 liste.append(i)             if i.R1 != None and i.R1 != "":         for i in listedossiers:     if (ch=="R1"):     listedossiers =DosTAff()     liste=[]          ch=request.GET.get('reg') def filtre_regT(request):            return render(request,"dossieratrait.html",context)          context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD}          NBD=nbrDAT()         veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(liste,9)                  liste.append(i)             if i.R14 != None and i.R14 != "":         for i in listedossiers:     elif (ch =="R14"):                                   liste.append(i)             if i.R13 != None and "doute rejeté" in i.R13 :         for i in listedossiers:     elif (ch =="R13_rejete"):                  liste.append(i)             if i.R13 != None and "doute confirmé" in i.R13 :         for i in listedossiers:     elif (ch =="R13_confirme"):                    liste.append(i)             if i.R12 != None and i.R12 != "":         for i in listedossiers:     elif (ch =="R12"):                 liste.append(i)             if i.R11 != None and i.R11 != "":         for i in listedossiers:     elif (ch =="R11"):                 liste.append(i)             if i.R10 != None and i.R10 != "":         for i in listedossiers:     elif (ch =="R10"):                 liste.append(i)             if i.R9 != None and i.R9 != "":         for i in listedossiers:     elif (ch =="R9"):                 liste.append(i)             if i.R8 != None and i.R8 != "":         for i in listedossiers:     elif (ch =="R8"):                 liste.append(i)             if i.R7 != None and i.R7 != "":         for i in listedossiers:     elif (ch =="R7"):                 liste.append(i)             if i.R6 != None and i.R6 != "":         for i in listedossiers:     elif (ch =="R6"):                 liste.append(i)             if i.R5 != None and i.R5 != "":         for i in listedossiers:     elif (ch =="R5"):                 liste.append(i) ad     �     Z       �  �  �  �  c  '      �  �  �  �  p  M  *    �  {  v  ?  >  =  <  ;  :  9  8  �  R  �  m  l  k  j  i  �
  ~
  
  �	  �	  �	  �	  �	  �	  ~	  {	  x	  u	  r	  q	  ^	  T	  	  �  �  }  Z     �  t  e  d  R  +  �  �  �  q  N  �  "    �  �  �  �  �  �  :  "  
     �  �  �  �  6     �  �  �                                              if (i.Statut!= "Changement procédure") and (i.RateFraude not in [0,0.0,None]):             i.RateFraude = str_to_float(i.RateFraude)             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:     Rate=0     list_veotest=veotest.objects.all()     NBD=0     list_Veo_recente=[]     NBDAT=test_nbrDAT()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def test_inis(request): @login_required       return NBD                 NBD=NBD+1             if ((Today_DateVeo-Date_création).days<=10 and (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté")   and i.Statut!="Dossier sans suite" and i.Statut!="Changement de procédure") :             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:     NBD=0     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_veotest=veotest.objects.all() def test_nbrDT():      return NBD                 NBD=NBD+1             if (((Today_DateVeo-Date_création).days<=5) and i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) :             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:     list_veotest=veotest.objects.all()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     NBD=0 def test_nbrDAT():  #  #  #  #  #  #  #  #  #  # * ####################################################################################################################" #####################################################################################################################* #################################################################################################################*#* ####################################################################################################################*     ################################################################################################################# ################################################################################################################## ################################################################################################################## ##################################################################################################################            return render(request,"dossiertrait.html",context)          context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBDAT}     NBDAT=nbrDAT()         veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(liste,9)                 liste.append(i)             if i.R14 != None and i.R14 != "":         for i in listedossiers:     elif (ch =="R14"):                                   liste.append(i)             if i.R13 != None and "doute rejeté" in i.R13 :         for i in listedossiers:     elif (ch =="R13_rejete"):                  liste.append(i)             if i.R13 != None and "doute confirmé" in i.R13 : ad  G   �     `       �  �  �  [  8    �  |  H  G  7    �  �  �  �  �  z  c  b  M  4        �  �  �  �  �  �  �  y  5        �  �  �  �  v  _  H  G  2         �
  �
  �
  �
  �
  �
  �
  �
  o
  n
  W
  <
  ;
  '
  
  �	  �	  �	  �	  �  �  t  \  R    �  �  {  X  �  �  r  c  b  P  )  �  �  �  o  L  �       �  �  �  �                                                                         def test_DosAff():      return NBD                 NBD=NBD+1             if ((Today_DateVeo-Date_création).days<=10 and (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté")   and i.Statut!="Dossier sans suite" and i.Statut!="Changement de procédure") :             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:     NBD=0     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_veotest=veotest.objects.all() def test_nbrDT():      return NBD                 NBD=NBD+1             if (((Today_DateVeo-Date_création).days<=5) and i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) :             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:     list_veotest=veotest.objects.all()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     NBD=0 def test_test_nbrDAT():     return render(request,"detail_test.html",context)      context={"SupUse":SupUse, "NBDT":NBDT,"NBDossiers":NBD,"Veo":Veo,"Rate":Rate ,"R1": R1,"R1_P": R1_P, "R1_A":R1_A, "R2":R2, "R2_DDA":R2_DDA, "R2_DS":R2_DS,"R3":R3, "R3_DDA":R3_DDA, "R3_DS":R3_DS, "R4":R4, "R4_SP":R4_SP, "R4_SA":R4_SA,"R5":R5 ,"R5_Assis":R5_Assis ,"R6":R6,"R6_Assis1":R6_Assis1 ,"R6_Assis2":R6_Assis2,"R7":R7,"R7_P":R7_P,"R7_A":R7_A, "R9_DFP":R9_DFP, "R9_DS":R9_DS, "R9":R9,"R8":R8,"R11":R11, "R10_Dos":R10_Dos,"R10":R10 , "R12_Dos":R12_Dos,"R12":R12 ,"R14":R14, "R13_Dos":R13_Dos,"R13":R13 }         SupUse = False     else:         SupUse = True     if request.user.is_superuser:     # Vérifier si c'est superuser     R14=Veo.Reg14()      R13_Dos=Veo.Reg13()[1]     R13=Veo.Reg13()[0]      R11=Veo.Reg11()      R12_Dos=Veo.Reg12()[1]     R12=Veo.Reg12()[0]          R10_Dos=Veo.Reg10()[1]     R10=Veo.Reg10()[0]      R8=Veo.Reg8()      R9_DS=Veo.Reg9()[2]     R9_DFP=Veo.Reg9()[1]     R9=Veo.Reg9()[0]      R7_A=Veo.Reg7()[2]     R7_P=Veo.Reg7()[1]     R7=Veo.Reg7()[0]      R6_Assis2=Veo.Reg6()[2]     R6_Assis1=Veo.Reg6()[1]     #Les  deux dossiers Assistance qui ne dépassent pas 3 mois     R6=Veo.Reg6()[0]      R5_Assis=Veo.Reg5()[1]     #Dossier assistance qui à la  date moins  de 7h et plus de 20h     R5=Veo.Reg5()[0]      R4_SA=Veo.Reg4()[2]     R4_SP=Veo.Reg4()[1]     R4=Veo.Reg4()[0]      R3_DS=Veo.Reg3()[2]     R3_DDA=Veo.Reg3()[1]     R3=Veo.Reg3()[0]      R2_DS=Veo.Reg2()[2]     R2_DDA=Veo.Reg2()[1]     R2=Veo.Reg2()[0]      R1_A=Veo.Reg1()[2]     R1_P=Veo.Reg1()[1]     R1=Veo.Reg1()[0]     NBDT=nbrDT()     NBD=test_nbrDAT()     Rate=Veo.RateFraude     Veo=get_object_or_404(veotest,id=Dossier) def test_details(request, Dossier): @login_required      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBDAT}     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                          list_Veo_recente.append(i) ad     }     U       �  l  T  -  ,    �  �  t  I  ,  +    �  �  m  F  E  *    �  x
  M
  0
  /
  
  �	  �	  �	  �	  v	  O	  2	  	  �  �  �  �  �  D  $  �  �  �  y  2    �  �  �    �  �  �  i  S  I  2         �  �  �  �  R  /  
     �  d  c  H  %    �  �  �  d  ?  5  �  �  �  }  |               def test_TrDsin(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=2     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrImmat(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg ,"tri":tri}     tri=1     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrDos(request):      return SupUse         SupUse = False     else:         SupUse = True     if request.user.is_superuser: def test_SupUse(request):     # Vérifier  si  l'utilisateur  connecter  est  un  admin     return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": list_Veo_recente}     #veopg.sort(key=lambda r: r.RateFraude,reverse=True)    # veopg = paginator.get_page(page)    # page = request.GET.get('page')    # paginator = Paginator(list_Veo_recente,9)         list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)             i.RateFraude=str_to_float(i.RateFraude)         for i in list_Veo_recente:     else:         list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     elif (id=="Date_sinistre"):         list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     if (id=="Date_creation"):     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff()     id=request.GET.get('filtre') def test_filtre(request):     return  list_Veo_recente             list_Veo_recente.append(i)         if i.statutdoute == "Doute confirmé":     for i in list_veotest:     NBD=test_nbrDAT()     list_veotest = veotest.objects.all()     list_Veo_recente =[] def test_DosAffdout():      return  list_Veo_recente                 list_Veo_recente.append(i)             if ((((Today_DateVeo-Date_création).days<=5) and (i.Statut!= "Changement procédure")) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" ) )and i.RateFraude not in [0,"0.0","","'0.0'",0.0,0,'0.0',None,'5.0','10.0']:             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:      list_veotest=veotest.objects.all()     list_Veo_recente=[]     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def test_DosAT():      return  list_Veo_recente                 list_Veo_recente.append(i)             if ((((Today_DateVeo-Date_création).days<=5) and (i.Statut!= "Changement procédure")) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" ) )and i.RateFraude not in [0,"0.0","","'0.0'",0.0,None]:             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:      list_veotest=veotest.objects.all()     list_Veo_recente=[]     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') ad  -   �     _       �  �  �  o  A    �  �  �  R  Q  8    �  �  �  x  U  0  &  �  �  �  n  K  5  $  �  �  �  j  `  �
  �
  �
  �
  �
  o
  ^
  
  �	  �	  �	  �	  5	  	   	  �  �  �  �  ]  /    �  �  t  @  ?  %    �  �  �  ^  ;      �  o  n  V  3      �  �  z  L  )    �  �  ]  \  =      �  �  �  ^  9  .  �  �                                                   context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=10     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrStatDoute(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=9     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrRF(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=8     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrIAdv(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=7     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrExp(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=6     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrStat(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=5     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrType(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=4     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrDcr(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=3     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() ad  .   �     a       �  �  �  �  y  h  $  �  �  �  �  9        �  �  �  �  d  6    �  �  {  G  F  *    �  �  �  j  G  "    �
  z
  y
  ^
  ;
  %
  
  �	  �	  }	  X	  M	  �  �  �  �  r  \  K    �  �  �  �    �  �  �  �  �  �  =    �  �  �  S        �  �  �  z  L  )    �  �  \  [  A      �  �  �  g  B  7  �  �                                                    context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=18     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrExpI(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=17     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrStatI(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=16     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrTypeI(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrDcrI(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrDsinI(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=13     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrImmatI(request):      return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg, "tri":tri}     tri=12     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrDosI(request):       return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg , "tri":tri}     tri=11     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_Trobs(request):      return render(request,"home_test.html",context) ad      �     ^       �  �  �  �  w  f    �  �  �  �  ,  �  �  �  �  �  v  F    �  �  �  �    �  �  �  �  z  5    �
  �
  �
  K
  
  �	  �	  �	  �	  n	  @	  	  �  �  �  P  O  N  M  2    �  �  �    \  7  -  �  �  �  j  H  2  !  �  �  �  b  X  �  �  �  t  ^  M    �  �  �  �    �  �  �  �  |  4    �  �  �  �                                      tri=4     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrDcrAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=3     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrDsinAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=2     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrImmatAT(request):      return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg ,"tri":tri}     tri=1     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrDosAT(request):        return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=22     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrobsI(request):     return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=21     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrStatDouteI(request):     return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=20     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=False)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrRFI(request):     return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=19     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAff() def test_TrIAdvI(request):      return render(request,"home_test.html",context) ad  /   �     [       �  Z  Y  =      �  �  �  _  :  0  �  �  n  L  6  %  �  �  �  o  e  �  �  �  �  l  [    �
  �
  �
  �
  2
  �	  �	  �	  �	  �	  �	  @	  	  �  �  �  W       �  �  �  �  h  %  �  �  �  �  <  �  �  �  �  �  Q  #     �  �  g  *      �  �  �  �  S  0       �  Y  X  W  ;      �  �  �                                                     list_Veo_recente.sort(key=lambda r: r.id,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrDosIAT(request):       return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg , "tri":tri}     tri=11     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT()  def test_TrobsAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=10     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrStatDouteAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=9     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrRFAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=8     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrIAdvAT(request):      return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=7     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrExpAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=6     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrStatAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=5     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrTypeAT(request):      return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri} ad     �     [       �  �  �      �  �  �  �  �  r  *  �  �  �  �  @    �  �  �  �  W  )    �  �  m  0  /    �
  �
  �
  �
  U
  2
  
  
  �	  \	  ?	  	  	  �  �  �  b  =  2  �  �  o  M  7  &  �  �  �  q  f  �  �  �  �  l  [    �  �  �  �  2  �  �  �  �  �  �  >    �  �  �  T    �  �  �  �  �  �                  for i in list_Veo_recente:     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrRFIAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=19     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrIAdvIAT(request):      return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=18     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrExpIAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=17     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrStatIAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=16     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrTypeIAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrDcrIAT(request):      return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrDsinIAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=13     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=True)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrImmatIAT(request):      return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg, "tri":tri}     tri=12     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9) ad  (   �     [       �  �  ^  ;      �  n  L  G  %    �  �  �  h  C  8  �  �  �  `  J  9  �  �  �  ~  s  �
  �
  �
  �
  �
  �
  k
  Z
  
  �	  �	  �	  �	  y	  b	  I	  	  �  �  �  b  =  �  t  s  W  3      �  �  r  M  C      �  �  �  Y  ,    �  U    �  �  �  �  l  >    �  �  �  �  �  h  C    �  �  �                                              pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=3     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDsinT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=2     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrImmatT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=1     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDosT(request):       return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri,"NBDT":NBDT}     tri=22     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT() def test_TrobsIAT(request):     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=21     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=False)     NBDT=nbrDT()     nbr=test_nbrDAT()     list_Veo_recente=test_DosAT()      def test_TrStatDouteIAT(request):     return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=20     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=False)         i.RateFraude=str_to_float(i.RateFraude) ad  
   �     X       �  N    �  �  �  �  e  7    �  �  �  �  �  a  <  �  �  �  �  �  �  �  �  {  e  T    �
  �
  �
  �
  k
  T
  ;
  
  �	  �	  y	  T	  /	  �  f  e  J  &    �  �  �  n  I  ?      �  �  �  U  (    �  Q    �  �  �  �  p  B    �  �  �  �  �  l  G    �  �  �    �  �  �  �  �                list_Veo_recente=test_DosTAff() def test_TrIAdvT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=7     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrExpT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=6     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrStatT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=5     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrTypeT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=4     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDcrT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD) ad     �     [       �  �  �  \  9    
  �  �  �  �  a     �  �  �    �  �  �  �  |  ]  -  �  �  �  t  j  E  .    �
  �
  �
  S
  .
  	
  |	  @	  ?	  	  �  �  �  �  b  ?      �  �  �  �  f  %  �  �  �  !  �  �  �  �  �    ;    �  �  �  �  ~  e  6    �  �  ~  Y  �  �  �  �  s  O  9  (  �  �  �  �                          page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDosIT(request):       return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=11     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff()  def test_TrobsT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=10     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrStatDouteT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=9     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrRFT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=8     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT() ad  =   �     Z       �  �  �  �  {  L  '  �  �  �  o  �  �  �  �  d  N  =  �  �  �    t  O  8    �  �  �  ]  8    �
  J
  .
  

  �	  �	  �	  o	  L	  '	  	  �  �  �  �  s  2    �  �  .  �  �  �  �  �  �  D    �  �  �  �  �  n  ?    �  �  �  b  �  �  �  |  X  B  1  �  �  �  u  j  E  .    �  �  �                                                                           list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDsinIT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDcrIT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDsinIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=13     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrImmatIT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=12     veopg = paginator.get_page(page) ad  �   �     U       �  �  m  H  �    ~  c  ?  )    �  �  �  [  P  +    �  �  �  f  9    �  b  &  
  �
  �
  �
  |
  N
  +
  
  �	  �	  �	  �	  w	  R	  	  �  �  �    �  �  �  {  j  +  �  �  �  �  �  n  U  &    �  �  n  I  �  �  e  A  +    �  �  �  e  Z  5      �  �  p  C    �  �                                                                                                                                               veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=18     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrExpIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=17     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrStatIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=16     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrTypeIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrDcrIT(request):      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True) ad     v     V       s  7    �  �  �  �  R  /  
  �  �  �  �  {  V    �  �  �    �  �  �  �  p  Q  !  �
  �
  �
  �
  ^
  S
  .
  
  �	  �	  �	  i	  <	  	  �  e  )    �  �  �  x  J  '    �  �  �  �  s  N    �  �  �  	  �  �  �  x  g  "  �  �  �  �  |  e  L    �  �  �  e  @  �  w  v             return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=22     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrobsIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=21     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrStatDouteIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=20     veopg = paginator.get_page(page)     page = request.GET.get('page')              paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=False)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrRFIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=19     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrIAdvIT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri} ad     �     Y       �  �  �  �  V  (    �  �  �  �  �  Q  ,  �  �  �  t  �  �  �  l  V  E    �  �  �  �  ]  F  -  �
  �
  �
  k
  F
  !
  �	  X	  H	  +	  	  �    i  X  :    �  �  q  \  E  0  &  
  �  �  z  �  �  �  @    �  �  �  k  7  '    �  �  \  F  5    �  �  [  B  )    �  �  �  �  �  �                      if i.Date_création!=None:         for i in liste:             liste=liste1+liste2         else:             liste=liste1         elif liste2==None:             liste=liste2         if liste1==None:         liste1=list(veotest.objects.filter(Immatriculation__icontains=query))         liste2=list(veotest.objects.filter(Dossier__icontains=query))         query=request.GET.get('search')     if request.method=='GET':     NBDT=nbrDT()     NBD=test_nbrDAT()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_Veo_recente=[] def test_filterDosAT(request): @login_required     return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD,"NBDT":NBDT}      veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                 i.RateFraude=str_to_float(i.RateFraude)                 list_Veo_recente.append(i)             if ((Today_DateVeo-Date_création).days<=100) and i.RateFraude not in [0,'0.0',None,'5.0','10.0','15.0'] and i not in list_Veo_recente:             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in liste:         liste=liste1+liste2     else:         liste=liste1     elif liste2==None:         liste=liste2     if liste1==None:     liste1=list(veotest.objects.filter(Immatriculation__icontains=query))     liste2=list(veotest.objects.filter(Dossier__icontains=query))         query=request.GET.get('search')     if request.method=='GET':     NBDT=nbrDT()     NBD=test_nbrDAT()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_Veo_recente=[] def test_filterDos(request): @login_required     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=23     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r:  r.date_obs,reverse=True)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrdateT(request):     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()     tri=24     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r:  r.date_obs,reverse=False)     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=test_DosTAff() def test_TrdateIT(request): ad     O     K       �  d  �  �  �  D    �  �  p  3  #    �  �  �    2    �
  �
  X
  ?
  &
  
  �	  �	  �	  �	  �	  (	  �  �  �  z  7  	  �  �  �  �  �    f  7    �  �    Z  �  �  �  �  j  T  C  +    �  �  ,  �  �  �  �  ]  :      �  �  �  �  O  N             list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]      veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)              list_Veo_recente.append(i)             i.RateFraude = str_to_float(i.RateFraude)         if (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté") and i.Statut!="Changement de procédure" and  i.Statut!="Dossier sans suite" :     for i in list_veotest:     Veoservice=veotest.objects.all()     list_veotest=test_DosTAff()     list_Veo_recente=[]     NBDT=nbrDT()     NBD=test_nbrDAT() def test_dossierstrait(request): @login_required      return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=veotest.objects.all()           veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                         i.RateFraude=str_to_float(i.RateFraude)                         list_Veo_recente.append(i)                     if (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté") and i.Statut!="Changement de procédure" and  i.Statut!="Dossier sans suite" and i.RateFraude not in [0,'0.0',None,'5.0','10.0'] and i not in list_Veo_recente:                 if ((Today_DateVeo-Date_création).days<=100):                 Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')             if i.Date_création!=None:         for i in liste:             liste=liste1+liste2         else:             liste=liste1         elif liste2==None:             liste=liste2         if liste1==None:         liste1=list(veotest.objects.filter(Immatriculation__icontains=query))         liste2=list(veotest.objects.filter(Dossier__icontains=query))         query=request.GET.get('search')     if request.method=='GET':     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     NBDT=nbrDT()     NBD=test_nbrDAT()     list_Veo_recente=[] def test_filterDosT(request): @login_required     return render(request,"dossieratrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD,"NBDT":NBDT}     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                         i.RateFraude=str_to_float(i.RateFraude)                         list_Veo_recente.append(i)                     if (i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) and i not in list_Veo_recente:                 if ((Today_DateVeo-Date_création).days<=100):                 Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M') ad     �     U       �  �  �    �  �  �  �  r  Z  I  *  �  �  �  |  a  X    �  �  �  �  u  G  $  �
  �
  P
  
  
  �	  �	  i	  Q	  *	  )	  	  �  �  �  �  �    X  /  �  �  �  W  
  �  �  �  �  r  X    �  �  �  @  6  �  �  �  g  E  /  �  �  �  �  s  \  [  6        �  �  �  �  �  �                              R4=round((Veo.Reg4()[0]*3)/15,2)      R3_DS=Veo.Reg3()[2]     R3_DDA=Veo.Reg3()[1]     R3=round((Veo.Reg3()[0]*2)/15,2)      R2_DS=Veo.Reg2()[2]     R2_DDA=Veo.Reg2()[1]     R2=round((Veo.Reg2()[0]*2)/15,2)      R1_A=Veo.Reg1()[2]     R1_P=Veo.Reg1()[1]     R1=round((Veo.Reg1()[0]*3/15),2)     Rate=Veo.RateFraude     Veo=get_object_or_404(veotest,id=dos)         veotest.objects.filter(id=dos).update(date_obs=dateM)        #dateM = ls[1]         #ls=str(dateM).split('.')         dateM=datetime.datetime.now()         veotest.objects.filter(id=dos).update(observation=query)     if query not in [None,""]:         veotest.objects.filter(id=dos).update(statutdoute="Non traité")     else:         veotest.objects.filter(id=dos).update(statutdoute="Pas sur")     elif (obs=="Pas sur"):         veotest.objects.filter(id=dos).update(statutdoute="Attente photos Avant")     elif (obs=="Attente"):         veotest.objects.filter(id=dos).update(statutdoute="Doute rejeté")     elif (obs=="rejete"):         veotest.objects.filter(id=dos).update(statutdoute="Doute confirmé")     if (obs=="confirme"):     ls=[]     NBDT=nbrDT()     NBD=test_nbrDAT()     veotest.objects.filter(id=dos).update(email_traitement=email_traitement)     veotest.objects.filter(id=dos).update(utilisateur=utilisateur)     dos=request.GET.get('dos')     email_traitement=request.user.username.title     utilisateur=request.user.first_name +" "+ request.user.last_name     query=request.GET.get('observation')     obs=request.GET.get('statutdoute') def test_observation(request):     return  list_Veo_recente                 list_Veo_recente.append(i)             if ((Today_DateVeo-Date_création).days<=8) and (i.Statut!= "Changement procédure") and  (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté"):             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_veotest:      list_veotest=veotest.objects.all()     list_Veo_recente=[]     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def test_DosTAff():      return render(request,"dossieratrait_test.html",context)      context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD,"NBDT":NBDT ,"list_inst": list_inst}    # veopg.sort(key=lambda r: r.RateFraude,reverse=True)     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)               list_Veo_recente.append(i)             i.RateFraude = str_to_float(i.RateFraude)         if (i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) :              for i in list_veotest:             list_inst.append(i)         if i.Statut =="Dossier en instruction" and "D" in i.Dossier:     for i in list_veotestall:     list_veotestall= veotest.objects.all()     list_veotest=test_DosAff()     list_inst=[]     list_Veo_recente=[]     NBDT=nbrDT()     NBD=test_nbrDAT() def test_dossiersAtrait(request): @login_required     return render(request,"dossiertrait_test.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9) ad  
        x       �  �  �  �  �  �  i  M  1  0      �  �  �  �  �  �  �  �  �  z  _  Z  C  (  '      �  �  �  �  �  �  �  �  �  m  O  J  =    	  �
  �
  �
  �
  g
  ;
  
  
  �	  �	  �	  �	  z	  Z	  .	  	  �  �  �  �  v  V  *  
  �  �  �  �  r  R  &    �  �  �  �  m  M    �  �  �  �  z  c  C    �  �  �  �  r  R  Q  3    �  �  �  �  �  n  @     �  �  �  �  D                                          return render(request,"home_test.html",context)     context={"SupUse":SupUse(request),"NBDossiers":NBDAT,"list_Veo_recente": veopg }     NBDAT=test_nbrDAT()         veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(liste,9)                 liste.append(i)             if i.R14 != None and i.R14 != "":         for i in listedossiers:     elif (ch =="R14"):                                   liste.append(i)             if i.R13 != None and "doute rejeté" in i.R13 :         for i in listedossiers:     elif (ch =="R13_rejete"):                  liste.append(i)             if i.R13 != None and "doute confirmé" in i.R13 :         for i in listedossiers:     elif (ch =="R13_confirme"):                      liste.append(i)             if i.R12 != None and i.R12 != "":         for i in listedossiers:     elif (ch =="R12"):                 liste.append(i)             if i.R11 != None and i.R11 != "":         for i in listedossiers:     elif (ch =="R11"):                 liste.append(i)             if i.R10 != None and i.R10 != "":         for i in listedossiers:     elif (ch =="R10"):                 liste.append(i)             if i.R9 != None and i.R9 != "":         for i in listedossiers:     elif (ch =="R9"):                 liste.append(i)             if i.R8 != None and i.R8 != "":         for i in listedossiers:     elif (ch =="R8"):                 liste.append(i)             if i.R7 != None and i.R7 != "":         for i in listedossiers:     elif (ch =="R7"):                 liste.append(i)             if i.R6 != None and i.R6 != "":         for i in listedossiers:     elif (ch =="R6"):                 liste.append(i)             if i.R5 != None and i.R5 != "":         for i in listedossiers:     elif (ch =="R5"):                 liste.append(i)             if i.R4 != None and i.R4 != "":         for i in listedossiers:     elif (ch =="R4"):                          liste.append(i)             if i.R3 != None and i.R3 != "":         for i in listedossiers:     elif (ch =="R3"):                 liste.append(i)             if i.R2 != None and i.R2 != "":         for i in listedossiers:     elif (ch =="R2"):                 liste.append(i)             if i.R1 != None and i.R1 != "":         for i in listedossiers:     if (ch=="R1"):     listedossiers =test_DosAff()     liste=[]          ch=request.GET.get('reg') def test_filtre_reg(request):       return render(request,"detail_test.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"Veo":Veo,"Rate":Rate ,"R1": R1,"R1_P": R1_P, "R1_A":R1_A, "R2":R2, "R2_DDA":R2_DDA, "R2_DS":R2_DS,"R3":R3, "R3_DDA":R3_DDA, "R3_DS":R3_DS, "R4":R4, "R4_SP":R4_SP, "R4_SA":R4_SA,"R5":R5 ,"R5_Assis":R5_Assis ,"R6":R6,"R6_Assis1":R6_Assis1 ,"R6_Assis2":R6_Assis2,"R7":R7,"R7_P":R7_P,"R7_A":R7_A, "R9_DFP":R9_DFP, "R9_DS":R9_DS, "R9":R9,"R8":R8,"NBDossiers":NBD,"R11":R11, "R10_Dos":R10_Dos,"R10":R10 , "R12_Dos":R12_Dos,"R12":R12,"R14":R14, "R13_Dos":R13_Dos,"R13":R13 }      R14=Veo.Reg14()      R13_Dos=Veo.Reg13()[1]     R13=Veo.Reg13()[0]      R11=Veo.Reg11()      R12_Dos=Veo.Reg12()[1]     R12=Veo.Reg12()[0]          R10_Dos=Veo.Reg10()[1]     R10=Veo.Reg10()[0]      R8=Veo.Reg8()       R9_DS=Veo.Reg9()[2]     R9_DFP=Veo.Reg9()[1]     R9=Veo.Reg9()[0]      R7_A=Veo.Reg7()[2]     R7_P=Veo.Reg7()[1]     R7=Veo.Reg7()[0]      R6_Assis2=Veo.Reg6()[2]     R6_Assis1=Veo.Reg6()[1]     R6=round((Veo.Reg6()[0]*2)/15,2)      R5_Assis=Veo.Reg5()[1]     R5=round((Veo.Reg5()[0]*2)/15,2)      R4_SA=Veo.Reg4()[2]     R4_SP=Veo.Reg4()[1] ad     	     w       �  �  �  �  �  }  ]  1    �  �  �  �  y  Y  -      �  �  �  �  l  L        �  �  �  ~  h  H    �  �  �  �  z  d  D    �
  �
  �
  �
  s
  \
  <
  
  �	  �	  �	  �	  i	  f	  F	  &	  �  �  �  �  �  M  -  ,      �  �  �  �  r  O  *      �  �  w  v  u  p  Q  3  .  !  �  �  �  �  �  j  J    �  �  �  �  |  s  ]  =    �  �  �  �  o  Y  9    �  �  �  �  k  U  5  	                                 if i.R8 != None and i.R8 != "":         for i in listedossiers:     elif (ch =="R8"):                 liste.append(i)             if i.R7 != None and i.R7 != "":         for i in listedossiers:     elif (ch =="R7"):                 liste.append(i)             if i.R6 != None and i.R6 != "":         for i in listedossiers:     elif (ch =="R6"):                 liste.append(i)             if i.R5 != None and i.R5 != "":         for i in listedossiers:     elif (ch =="R5"):                 liste.append(i)             if i.R4 != None and i.R4 != "":         for i in listedossiers:     elif (ch =="R4"):                          liste.append(i)             if i.R3 != None and i.R3 != "":         for i in listedossiers:     elif (ch =="R3"):                 liste.append(i)             if i.R2 != None and i.R2 != "":         for i in listedossiers:     elif (ch =="R2"):                 liste.append(i)             if i.R1 != None and i.R1 != "":         for i in listedossiers:     if (ch=="R1"):     listedossiers =test_DosTAff()     liste=[]          ch=request.GET.get('reg') def test_filtre_regT(request):            return render(request,"dossieratrait_test.html",context)          context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD}          NBD=test_nbrDAT()         veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(liste,9)                  liste.append(i)             if i.R14 != None and i.R14 != "":         for i in listedossiers:     elif (ch =="R14"):                                   liste.append(i)             if i.R13 != None and "doute rejeté" in i.R13 :         for i in listedossiers:     elif (ch =="R13_rejete"):                  liste.append(i)             if i.R13 != None and "doute confirmé" in i.R13 :         for i in listedossiers:     elif (ch =="R13_confirme"):                    liste.append(i)             if i.R12 != None and i.R12 != "":         for i in listedossiers:     elif (ch =="R12"):                 liste.append(i)             if i.R11 != None and i.R11 != "":         for i in listedossiers:     elif (ch =="R11"):                 liste.append(i)             if i.R10 != None and i.R10 != "":         for i in listedossiers:     elif (ch =="R10"):                 liste.append(i)             if i.R9 != None and i.R9 != "":         for i in listedossiers:     elif (ch =="R9"):                 liste.append(i)             if i.R8 != None and i.R8 != "":         for i in listedossiers:     elif (ch =="R8"):                 liste.append(i)             if i.R7 != None and i.R7 != "":         for i in listedossiers:     elif (ch =="R7"):                 liste.append(i)             if i.R6 != None and i.R6 != "":         for i in listedossiers:     elif (ch =="R6"):                 liste.append(i)             if i.R5 != None and i.R5 != "":         for i in listedossiers:     elif (ch =="R5"):                 liste.append(i)             if i.R4 != None and i.R4 != "":         for i in listedossiers:     elif (ch =="R4"):                          liste.append(i)             if i.R3 != None and i.R3 != "":         for i in listedossiers:     elif (ch =="R3"):                 liste.append(i)             if i.R2 != None and i.R2 != "":         for i in listedossiers:     elif (ch =="R2"):                 liste.append(i)             if i.R1 != None and i.R1 != "":         for i in listedossiers:     if (ch=="R1"):     listedossiers =test_DosAT()     liste=[]          ch=request.GET.get('reg') def test_filtre_regAT(request): ad  "   �     h       �  �  �  ~  ^  G  '  �  �  �  �  t  T  =    �  �  �  �  �  N  .  -    �  �  �  �  �  j  J    �  �  �  �  �  t  �
  �
  �
  �
  o
  n
  W
  /
  .
  -
  ,
  
  �	  �	  �	  �	  �	  �	  \	  D	  J  4      �  �  {  z  \  3  )      �  �  �  u  j  T  =  �  u  n  D  2    c  E  .  y  d  G  *    �  �  �  t  h  c  H  ?  )  �  �  �  �                                             response=ls     ls = serialize('json', Veoservices.objects.all())         #ls.append(i)              #for i in  veoservice:          #ls =[]     veoservice=Veoservices.objects.all() def  getVeos(request):     return HttpResponse(response, content_type='text/json')"""     response = jsls     #jsl = [line for line in jsls]     #jsls = json.loads(jsls)     #jsls = json.dumps(jsls)     jsls.append(']')     jsls.append({'Dossier':l.Dossier,'Pourcentage Fraude':l.RateFraude,'Procédure':l.Procédure,'Statut':l.Statut,'Date Création':l.Date_création,'Statut doute':l.statutdoute})      jsls.append(",")               jsls.append(js)               js={'Dossier':j.Dossier,'Pourcentage Fraude':j.RateFraude,'Procédure':j.Procédure,'Statut':j.Statut,'Date Création':j.Date_création,'Statut doute':j.statutdoute}             jsls.append(",")             N=N+1         if  j != k and j != l and N<1001:            for j  in  ls:     jsls.append({'Dossier':k.Dossier,'Pourcentage Fraude':k.RateFraude,'Procédure':k.Procédure,'Statut':k.Statut,'Date Création':k.Date_création,'Statut doute':k.statutdoute})      jsls.append('[')       l=ls[len(ls)-1]                  k=ls[0]             ls.append(i)         if i.RateFraude not in ["0.0",0.0,None,"0",0,"5.0",5.0,5,"10.0",10.0,10,"15.0",15.0,15]:     for i in  veoservice:     N=2     jsls=[]     ls=[]     veoservice=Veoservices.objects.all() """def get_dossiers(request):      return HttpResponse(response, content_type='text/json')     response = json.loads(response)                 response =  json.dumps([{'Error':Dossier}])              if veo == None:                 break                 response = json.dumps([{'Dossier':Dossier,'Immatriculation':veo.Immatriculation,'Pourcentage Fraude':veo.RateFraude,'Procédure':veo.Procédure,'Statut':veo.Statut,'Date Création':veo.Date_création,'Statut doute':veo.statutdoute}])                 veo = i             if i.Dossier == Dossier:         for i in  veoservice:                      if request.method == 'GET':     veo=None     veoservice=Veoservices.objects.all() def get_veoservices(request,Dossier):        return render(request,"index.html") def template(request):  ################## Affichage du  templates  ##############"##############"      return render(request,"dossiertrait_test.html",context)          context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": test_DosAffdout(),"NBDossiers":NBDAT}     NBDAT=test_nbrDAT()         veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(liste,9)                  liste.append(i)             if i.R14 != None and i.R14 != "":         for i in listedossiers:     elif (ch =="R14"):                                   liste.append(i)             if i.R13 != None and "doute rejeté" in i.R13 :         for i in listedossiers:     elif (ch =="R13_rejete"):                  liste.append(i)             if i.R13 != None and "doute confirmé" in i.R13 :         for i in listedossiers:     elif (ch =="R13_confirme"):                    liste.append(i)             if i.R12 != None and i.R12 != "":         for i in listedossiers:     elif (ch =="R12"):                 liste.append(i)             if i.R11 != None and i.R11 != "":         for i in listedossiers:     elif (ch =="R11"):                 liste.append(i)             if i.R10 != None and i.R10 != "":         for i in listedossiers:     elif (ch =="R10"):                 liste.append(i)             if i.R9 != None and i.R9 != "":         for i in listedossiers:     elif (ch =="R9"):                 liste.append(i) ad  3   �     b       �  �  �  �  (  �  �  �  f  Y    �  �  �  U    �  �  �  �  p  X  G  6  !  
  �  �  �  �  �  �  �  }  e  d  O  7      	  �
  �
  �
  �
  T
  8
  
  
  
  �	  �	  �	  �	  �	  �	  �	  ~	  }	  f	  K	  F	  /	  	  	  �  �  �  �  �  �  �  q  [  Q  :  :  9    �  �  �  [  ,    �  �      �  �  �  �  q  #    �  �  �                                                             if i.Date_création!=None:     for i in list_Veoservices:     NBD=0     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_Veoservices=Veoservices.objects.all() def nbrDT():      return NBD                 NBD=NBD+1             if (((Today_DateVeo-Date_création).days<=5) and i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) :             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_Veoservices:     list_Veoservices=Veoservices.objects.all()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo, '%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     NBD=0 def nbrDAT():     return render(request,"detail.html",context)      context={"SupUse":SupUse, "NBDT":NBDT,"NBDossiers":NBD,"Veo":Veo,"Rate":Rate ,"R1": R1,"R1_P": R1_P, "R1_A":R1_A, "R2":R2, "R2_DDA":R2_DDA, "R2_DS":R2_DS,"R3":R3, "R3_DDA":R3_DDA, "R3_DS":R3_DS, "R4":R4, "R4_SP":R4_SP, "R4_SA":R4_SA,"R5":R5 ,"R5_Assis":R5_Assis ,"R6":R6,"R6_Assis1":R6_Assis1 ,"R6_Assis2":R6_Assis2,"R7":R7,"R7_P":R7_P,"R7_A":R7_A, "R9_DFP":R9_DFP, "R9_DS":R9_DS, "R9":R9,"R8":R8,"R11":R11, "R10_Dos":R10_Dos,"R10":R10 , "R12_Dos":R12_Dos,"R12":R12 , "R13_Dos":R13_Dos,"R13":R13, "R14":R14}         SupUse = False     else:         SupUse = True     if request.user.is_superuser:     # Vérifier si c'est superuser     R14 =Veo.Reg14()      R13_Dos=Veo.Reg13()[1]     R13=Veo.Reg13()[0]      R11=Veo.Reg11()      R12_Dos=Veo.Reg12()[1]     R12=Veo.Reg12()[0]          R10_Dos=Veo.Reg10()[1]     R10=Veo.Reg10()[0]      R8=Veo.Reg8()      R9_DS=Veo.Reg9()[2]     R9_DFP=Veo.Reg9()[1]     R9=Veo.Reg9()[0]      R7_A=Veo.Reg7()[2]     R7_P=Veo.Reg7()[1]     R7=Veo.Reg7()[0]      R6_Assis2=Veo.Reg6()[2]     R6_Assis1=Veo.Reg6()[1]     #Les  deux dossiers Assistance qui ne dépassent pas 3 mois     R6=Veo.Reg6()[0]      R5_Assis=Veo.Reg5()[1]     #Dossier assistance qui à la  date moins  de 7h et plus de 20h     R5=Veo.Reg5()[0]      R4_SA=Veo.Reg4()[2]     R4_SP=Veo.Reg4()[1]     R4=Veo.Reg4()[0]      R3_DS=Veo.Reg3()[2]     R3_DDA=Veo.Reg3()[1]     R3=Veo.Reg3()[0]      R2_DS=Veo.Reg2()[2]     R2_DDA=Veo.Reg2()[1]     R2=Veo.Reg2()[0]      R1_A=Veo.Reg1()[2]     R1_P=Veo.Reg1()[1]     R1=Veo.Reg1()[0]     NBDT=nbrDT()     NBD=nbrDAT()     Rate=Veo.RateFraude     Veo=get_object_or_404(Veoservices,id=Dossier) def details(request, Dossier): @login_required      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBDAT}     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)                          list_Veo_recente.append(i)                      if (i.Statut!= "Changement procédure") and (i.RateFraude not in [0,0.0,None]):             i.RateFraude = str_to_float(i.RateFraude)             i.Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_Veoservices:     Rate=0     list_Veoservices=Veoservices.objects.all() ad     v     S       �  �  �  �  �  �  U    �  �  �  �  ~  %    �  �  �  �  f      �
  �
  �
  �
  6
  �  �  �  �  �  �  Z  I  *  �  �  �  �  �  c  R  A  #  �  �  n  d  A    �  �  s  M    �  |  >  )    �  �  �  �  �  �  �  z  i  -  �  �  �  �  E      �  �  �  �  v  u                    list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrImmat(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg ,"tri":tri}     tri=1     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrDos(request):      return SupUse         SupUse = False     else:         SupUse = True     if request.user.is_superuser: def SupUse(request):     # Vérifier  si  l'utilisateur  connecter  est  un  admin     return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": list_Veo_recente}     #veopg.sort(key=lambda r: r.RateFraude,reverse=True)    # veopg = paginator.get_page(page)    # page = request.GET.get('page')    # paginator = Paginator(list_Veo_recente,9)         list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)             i.RateFraude=str_to_float(i.RateFraude)         for i in list_Veo_recente:     else:         list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     elif (id=="Date_sinistre"):         list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     if (id=="Date_creation"):     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff()     id=request.GET.get('filtre') def filtre(request):     return  list_Veo_recente             list_Veo_recente.append(i)         if i.statutdoute == "Doute confirmé":     for i in list_Veoservices:     NBD=nbrDAT()     list_Veoservices = Veoservices.objects.all()     list_Veo_recente =[] def DosAffdout():      return  list_Veo_recente                 list_Veo_recente.append(i)             if ((((Today_DateVeo-Date_création).days<=25) and (i.Statut!= "Changement procédure")) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" ) )and i.RateFraude not in [0,"0.0","","'0.0'",0.0,0,'0.0',None,'5.0','10.0']:             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_Veoservices:      list_Veoservices=Veoservices.objects.all()     list_Veo_recente=[]     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def DosAT():      return  list_Veo_recente                 list_Veo_recente.append(i)             if ((((Today_DateVeo-Date_création).days<=10) and (i.Statut!= "Changement procédure")) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" ) )and i.RateFraude not in [0,"0.0","","'0.0'",0.0,None]:             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_Veoservices:      list_Veoservices=Veoservices.objects.all()     list_Veo_recente=[]     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def DosAff():      return NBD                 NBD=NBD+1             if ((Today_DateVeo-Date_création).days<=10 and (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté")   and i.Statut!="Dossier sans suite" and i.Statut!="Changement de procédure") :             Date_création=datetime.datetime.strptime(i.Date_création, '%d/%m/%Y %H:%M') ad     �     d       �  �  �  �    �  �  �  �  �  �  K    �  �  �  b  3  2       �  �  �  h  E       �  ~  }  h  J  9  (  �
  �
  �
  n
  d
  �	  �	  �	  �	  �	  �	  v	  6	  	  �  �  �  M      	  �  �  �  �  [  8    	  �  q  p  [  =  ,    �  �  {  V  L  �  �  �  �  �  q  `  A    �  �  }  X  N  �  �  �  �  }  l  [    �  �  �                                page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrStatDoute(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=9     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrRF(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=8     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrIAdv(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=7     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrExp(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=6     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrStat(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=5     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrType(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=4     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrDcr(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=3     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrDsin(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=2     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9) ad  )   �     d       �  �  g  8  7  #    �  �  �  q  N  )    �  �  �  �  n  P  ?  .  �  �  �  }  r  
  �  �  �  �  �  �  ;    �
  �
  �
  Q
  "
  !
  
  �	  �	  �	  �	  W	  4	  	  	  �  l  k  V  8  '    �  �  ~  Y  N  �  �  �  �  �  p  _    �  �  �  �  2      �  �  �  �  m  ?    �  �  �  T  S  >       �  �  �  n  I  >  �  �                                               context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=18     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrExpI(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=17     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrStatI(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=16     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrTypeI(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrDcrI(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrDsinI(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=13     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrImmatI(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg, "tri":tri}     tri=12     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrDosI(request):       return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg , "tri":tri}     tri=11     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def Trobs(request):      return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=10     veopg = paginator.get_page(page) ad     �     a       �  �  �  �  �  z  *  �  �  �  �  @    �  �  �  �  �  n  *  �  �  �  �  @    �  �  �  �  q  C     �
  �
  �
  X
  C
  %
  
  
  �	  �	  m	  H	  =	  �  �  �  �  �  �  o  ^  M    �  �  �  �  )  �  �  �  �  �  �  P  "  �  �  �  g  /    �  �  �  �  d  A      �  q  [  >  -    �  �  �  ^  T  �  �  �  �                         return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=4     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrDcrAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=3     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrDsinAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=2     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrImmatAT(request):      return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg ,"tri":tri}     tri=1     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrDosAT(request):        return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=22     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrobsI(request):     return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=21     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrStatDouteI(request):     return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=20     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=False)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrRFI(request):     return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=19     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAff() def TrIAdvI(request):      return render(request,"home.html",context) ad     �     a       �  �  �  �  f  8    �  �  }  E  .       �  �  �  ^  9  /  �  �  x  [  J  9  �  �  �  �  y    �
  �
  �
  �
  �
  �
  2
  
  �	  �	  �	  I	  	  �  �  �  �  �  n  +  �  �  �  �  B  
  �  �  �  �  k  =    �  �  �  I  3  2      �  �  �  ^  9  .  �  �  �  �  s  V  E  4  �  �  �  �  x    �  �  �  �           list_Veo_recente=DosAT() def TrImmatIAT(request):      return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente":veopg, "tri":tri}     tri=12     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrDosIAT(request):       return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg , "tri":tri}     tri=11     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT()  def TrobsAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=10     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrStatDouteAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=9     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrRFAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=8     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrIAdvAT(request):      return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=7     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrExpAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=6     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrStatAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=5     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrTypeAT(request): ad     �     _       �  �  �  h  E       �  t  \  ?  .    �  �  �  a  V  �  �  �  �  �  o  ^    �  �  �  �  -  �
  �
  �
  �
  �
  [
  -
  

  �	  �	  q	  9	  !	  	  �  �  �  u  R  -  "  �  �  j  M  <  +  �  �  �  v  k    �  �  �  �  �  r  "  �  �  �  �  8     �  �  �  �  �  \    �  �  �  �  .  �  �  �  �  �  �  �            NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT()      def TrStatDouteIAT(request):     return render(request,"home.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=20     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=False)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrRFIAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=19     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrIAdvIAT(request):      return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=18     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrExpIAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=17     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrStatIAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=16     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrTypeIAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrDcrIAT(request):      return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrDsinIAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=13     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=True)     NBDT=nbrDT()     nbr=nbrDAT() ad     �     ]       �  �  j  E  :  �  �  �  q  `  O  
  �  �  �  �    �  �  �  �  �  �  �  H    �  �  �  �  �  o  @    �
  �
  �
  c
  �	  �	  �	  �	  m	  \	  K	  	  �  �  �  �  Y  B  )  �  �  �  g  B    �  ^  H  )      �  �  o  J  @       �  �  �  R  %     �  S      �  �  �  ~  P  -    �  �  �  �  �                           for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=4     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDcrT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=3     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDsinT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=2     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrImmatT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=1     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDosT(request):       return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDT":NBDT,"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri,"NBDT":NBDT}     tri=22     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=False)     NBDT=nbrDT()     nbr=nbrDAT()     list_Veo_recente=DosAT() def TrobsIAT(request):     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"NBDossiers":nbr,"list_Veo_recente": veopg, "tri":tri}     tri=21     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=False) ad  s   �     Y       �  �  k  >    �  l  5  4    �  �  �  �  k  H  #    �  �  �  �  l  +  �  �  �  ,  �
  �
  �
  �
  �
  �
  ]
  /
  
  �	  �	  �	  �	  �	  U	  0	  �  �  �  x  �  �  �  �  t  c  #  �  �  �  �  z  c  J    �  �  �  c  >  �    ~  h  I  8  '  �  �  �  b  X  /    �  �  �  j  =    �  �                                                                                                                         veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=8     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrIAdvT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=7     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrExpT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=6     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrStatT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=5     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrTypeT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé": ad     �     ]       x  A  -    �  �  �  �  Z  ,  	  �  �  �  �  �  R  -  �  �  �  u  �  �  �  �  {  j  Y    �
  �
  �
  �
  k
  T
  ;
  
  �	  �	  y	  T	  /	  �  p  [  Z  ;  *    �  �  �  _  T  +    �  �  �  f  9    �  g  0  /  .    �  �  �  �  n  K  &    �  �  �  �  n  -     �  �  .  �  �  �  �  �  �  �                   NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrImmatIT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=12     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.id,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDosIT(request):       return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=11     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff()  def TrobsT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=10     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrStatDouteT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=9     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrRFT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri} ad     �     \       �  �  g  B  7    �  �  �  �  I    �  �  J    �  �  �  �  u  G  $  �  �  �  �  �  l  G    �
  �
  �
  
  �	  �	  �	  �	  �	  x	  1	  	  �  �  �  �  p  W  (    �  �  p  K  �  �  �  t  U  D  3  �  �  �  w  l  C  ,    �  �  ~  Q  ,      H  G  1      �  �  {  X  3  (  �  �  �  �  �                              if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDcrIT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDsinIT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=15     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_création,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDcrIT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=14     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Date_sinistre,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrDsinIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=13     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Immatriculation,reverse=True) ad  #   �     V       �  �  m  H  #  �  d  M  .      �  �  x  S  H      �  �  �  Z  -    �  [  $    �
  �
  �
  �
  _
  <
  
  
  �	  �	  �	  �	  _	  	  �  �  �    �  �  �  �  �  R  $    �  �  �  �  x  I  $  �  �  �  l  �  �  �  w  f  U    �  �  �  �  [  D  +  �  �  �  i  D    �  �                                         context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=19     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.ImmatriculationAdverse,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrIAdvIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=18     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Expert,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrExpIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=17     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Statut,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrStatIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=16     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.Procédure,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrTypeIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i) ad     �     [       �  �  �  �  s  T  $  �  �  �  �  a  V  -    �  �  �  h  ;    �  i  2    �  �  �  �  b  ?      �
  �
  �
  �
  b
  !
  �	  �	  �	  "	  �  �  �  �  �  O  !  �  �  �  �  �  u  F  !  �  �  �  i  �  �  �  �  s  b  Q    �  �  �  �  d  M  4    �  �  r  M  (  �  i  S  4  #    �  �  �                                paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r:  r.date_obs,reverse=True)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrdateT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=24     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r:  r.date_obs,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrdateIT(request):      return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=22     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.observation,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrobsIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=21     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.statutdoute,reverse=False)     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrStatDouteIT(request):     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=20     veopg = paginator.get_page(page)     page = request.GET.get('page')              paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=False)         i.RateFraude=str_to_float(i.RateFraude)     for i in list_Veo_recente:     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=DosTAff() def TrRFIT(request):     return render(request,"dossiertrait.html",context) ad  ?   �     O       �  �  �  �  m  T  %     �  �  m  H  �  �  y  a  I    �  �  �  u  M    �  �  �  x  c  Y  =  )    �
  
  �	  �	  s	  E	  "	  �  �  �  o  _  E  -  �  �  �  w  Y  1  �  �  |  c  H  /  !    �  �  e  &  �  �  I    �  �  �  2  �  �  �  �  �  �  �                                                                     NBDT=nbrDT()     NBD=nbrDAT()     list_Veo_recente=[] def filterDosT(request): @login_required     return render(request,"dossieratrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD,"NBDT":NBDT}     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                         i.RateFraude=str_to_float(i.RateFraude)                         list_Veo_recente.append(i)                     if (i.statutdoute=="Non traité" and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) or (i.statutdoute=="Attente photos Avant" and i.Photos_Avant!="" and i.Photos_Avant!=None and i.Statut!="Changement de procédure" and i.RateFraude not in [0,'0.0',None,'5.0','10.0']) and i not in list_Veo_recente:                 if ((Today_DateVeo-Date_création).days<=100):                 Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')             if i.Date_création!=None:         for i in liste:             liste=liste1+liste2         else:             liste=liste1         elif liste2==None:             liste=liste2         if liste1==None:         liste1=list(Veoservices.objects.filter(Immatriculation__icontains=query))         liste2=list(Veoservices.objects.filter(Dossier__icontains=query))         query=request.GET.get('search')     if request.method=='GET':     NBDT=nbrDT()     NBD=nbrDAT()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_Veo_recente=[] def filterDosAT(request): @login_required     return render(request,"home.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD,"NBDT":NBDT}      veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)                 i.RateFraude=str_to_float(i.RateFraude)                 list_Veo_recente.append(i)             if ((Today_DateVeo-Date_création).days<=100) and i.RateFraude not in [0,'0.0',None,'5.0','10.0','15.0'] and i not in list_Veo_recente:             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in liste:         liste=liste1+liste2     else:         liste=liste1     elif liste2==None:         liste=liste2     if liste1==None:     liste1=list(Veoservices.objects.filter(Immatriculation__icontains=query))     liste2=list(Veoservices.objects.filter(Dossier__icontains=query))         query=request.GET.get('search')     if request.method=='GET':     NBDT=nbrDT()     NBD=nbrDAT()     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M')     list_Veo_recente=[] def filterDos(request): @login_required     return render(request,"dossiertrait.html",context)     context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"list_Veo_Doute": DosAffdout(),"NBDossiers":NBD,"NBDT":NBDT, "tri":tri}     veoD = paginator.get_page(pageD)     pageD = request.GET.get('pageD')     paginatorD = Paginator(list_Veo_Doute,9)     list_Veo_Doute.sort(key=lambda r: r.RateFraude,reverse=True)             list_Veo_Doute.append(i)         if i.statutdoute == "Doute confirmé":     for i in Veoservice:     list_Veo_Doute =[]     Veoservice=Veoservices.objects.all()     tri=23     veopg = paginator.get_page(page)     page = request.GET.get('page') ad  �  M     d       �  �  �  �  f  C    �  �  k  2  1  "  �  �  v  G  F  '    �  �  �  �  �  v  M    �
  �
  q
   
  
  �	  �	  �	  �	  o	   	  	  �  �  K  A  �  �  �  j  H  2  �  �  �  �  n  W  V  1       �  �  �  �  �  �  k  S  R  -      �  �  �  �  �  �  p  o  Z  A  )  (  '      �  �  �  �  �  �  �  �  ~  c  b  N  M  L                                                                                                                                                                                                                                                                                                                                                                                                                                        R14=Veo.Reg14()      R13_Dos=Veo.Reg13()[1]     R13=Veo.Reg13()[0]      R11=Veo.Reg11()      R12_Dos=Veo.Reg12()[1]     R12=Veo.Reg12()[0]          R10_Dos=Veo.Reg10()[1]     R10=Veo.Reg10()[0]      R8=Veo.Reg8()       R9_DS=Veo.Reg9()[2]     R9_DFP=Veo.Reg9()[1]     R9=Veo.Reg9()[0]      R7_A=Veo.Reg7()[2]     R7_P=Veo.Reg7()[1]     R7=Veo.Reg7()[0]      R6_Assis2=Veo.Reg6()[2]     R6_Assis1=Veo.Reg6()[1]     R6=round((Veo.Reg6()[0]*2)/15,2)      R5_Assis=Veo.Reg5()[1]     R5=round((Veo.Reg5()[0]*2)/15,2)      R4_SA=Veo.Reg4()[2]     R4_SP=Veo.Reg4()[1]     R4=round((Veo.Reg4()[0]*3)/15,2)      R3_DS=Veo.Reg3()[2]     R3_DDA=Veo.Reg3()[1]     R3=round((Veo.Reg3()[0]*2)/15,2)      R2_DS=Veo.Reg2()[2]     R2_DDA=Veo.Reg2()[1]     R2=round((Veo.Reg2()[0]*2)/15,2)      R1_A=Veo.Reg1()[2]     R1_P=Veo.Reg1()[1]     R1=round((Veo.Reg1()[0]*3/15),2)     Rate=Veo.RateFraude     Veo=get_object_or_404(Veoservices,id=dos)         Veoservices.objects.filter(id=dos).update(date_obs=dateM)        #dateM = ls[1]         #ls=str(dateM).split('.')         dateM=datetime.datetime.now()         Veoservices.objects.filter(id=dos).update(observation=query)     if query not in [None,""]:         Veoservices.objects.filter(id=dos).update(statutdoute="Non traité")     else:         Veoservices.objects.filter(id=dos).update(statutdoute="Pas sur")     elif (obs=="Pas sur"):         Veoservices.objects.filter(id=dos).update(statutdoute="Attente photos Avant")     elif (obs=="Attente"):         Veoservices.objects.filter(id=dos).update(statutdoute="Doute rejeté")     elif (obs=="rejete"):         Veoservices.objects.filter(id=dos).update(statutdoute="Doute confirmé")     if (obs=="confirme"):     ls=[]     NBDT=nbrDT()     NBD=nbrDAT()     Veoservices.objects.filter(id=dos).update(email_traitement=email_traitement)     Veoservices.objects.filter(id=dos).update(utilisateur=utilisateur)     dos=request.GET.get('dos')     email_traitement=request.user.username.title     utilisateur=request.user.first_name +" "+ request.user.last_name     query=request.GET.get('observation')     obs=request.GET.get('statutdoute') def observation(request):     return  list_Veo_recente                 list_Veo_recente.append(i)             if ((Today_DateVeo-Date_création).days<=8) and (i.Statut!= "Changement procédure") and  (i.statutdoute=="Doute confirmé" or i.statutdoute=="Doute rejeté"):             Date_création=datetime.datetime.strptime(i.Date_création,'%d/%m/%Y %H:%M')         if i.Date_création!=None:     for i in list_Veoservices:      list_Veoservices=Veoservices.objects.all()     list_Veo_recente=[]     Today_DateVeo=datetime.datetime.strptime(Today_DateVeo,'%d/%m/%Y %H:%M')     Today_DateVeo=datetime.datetime.today().strftime('%d/%m/%Y %H:%M') def DosTAff():      return render(request,"dossieratrait.html",context)      context={"SupUse":SupUse(request),"list_Veo_recente": veopg,"NBDossiers":NBD,"NBDT":NBDT ,"list_inst": list_inst}        # veopg.sort(key=lambda r: r.RateFraude,reverse=True)     veopg = paginator.get_page(page)     page = request.GET.get('page')     paginator = Paginator(list_Veo_recente,9)     list_Veo_recente.sort(key=lambda r: r.RateFraude,reverse=True)               list_Veo_recente.append(i) 